`timescale 1ns / 1ps

module test_memory;

    // parameters
    parameter BRAM_WIDTH = 10;
    parameter DATA_WIDTH = 32;

    logic clk;
    logic [2:0] op;
    logic [31:0] ab;
    logic [31:0] result;
    logic done;





endmodule